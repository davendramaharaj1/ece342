module part3
(
    input                       clk,
    input				        reset
);

endmodule
